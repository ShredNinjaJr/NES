
module pll (
	reset_reset_n,
	clk_clk,
	ppu_clk_clk,
	cpu_clk_clk,
	master_clk_clk);	

	input		reset_reset_n;
	input		clk_clk;
	output		ppu_clk_clk;
	output		cpu_clk_clk;
	output		master_clk_clk;
endmodule
