/* module that contains the CHR_ROM of the cartridge */
module CHR_ROM(clk, addr,data_out);
parameter n = 13;
parameter w = 8;

input clk;
input [n-1:0] addr;
output logic[w-1:0] data_out;

// Start module here!
reg [w-1:0] reg_array [2**n-1:0];
initial
begin
    $readmemh("../ROMs/dk_chr.txt", reg_array);
end



    assign data_out= reg_array[addr];
endmodule
